library verilog;
use verilog.vl_types.all;
entity muxTestBench is
end muxTestBench;
